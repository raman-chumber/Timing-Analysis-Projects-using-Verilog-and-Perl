`timescale 1ns/1ns
`include "d_ff.v";
`include "memory.v";

module memory_fixture;
reg [2:0] i;
reg [1:0] a;
reg cs, rd, oe;
wire [2:0] op;

reg [2:0] o;
reg [7:0] read [0:23];
reg [7:0] write [0:23];
integer m,j;

// Instantiate module 
memory m1(.cs(cs), .rd(rd), .oe(oe), .I(i), .A(a), .O(op));

// TASK 
task file_data;
input [7:0] read;
input [7:0] write;
 begin
  cs = write[7];
  oe = write[6];
  rd = write[5];
   a = {write[4],write[3]};
   i = {write[0],write[1],write[2]};
   #40;
  $display("WRITE op: cs=%b, oe=%b, rd=%b, a1=%b, a0=%b, i0=%b, i1=%b, i2=%b",cs,oe,rd,a[1],a[0],i[0],i[1],i[2]);
   #40;
  cs = read[7];
  oe = read[6];
  rd = read[5];
   a = {read[4],read[3]};
   o = {read[0],read[1],read[2]};
    #10;
  $display(" READ op: cs=%b, oe=%b, rd=%b, a1=%b, a0=%b, o0=%b, o1=%b, o2=%b",cs,oe,rd,a[1],a[0],op[0],op[1],op[2]);
 end
endtask

// MAIN
initial
 begin
 $readmemb("mem_op.txt",write); // Read from data file generated by Perl code
 $readmemb("mem_ip.txt",read);
 #40;

 for (j=0; j<=22; j=j+1)
  begin
   file_data(write[j],read[j]);
   #20;
   if (op === o)
      $display("Perl=%b: PASS\n",o);
   else
      $display("Perl=%b: FAIL\n",o);
  end
 end

initial
   #3000 $finish;
endmodule
